library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

package microcode_pkg is

type rom_t is array (0 to 2047) of STD_LOGIC_VECTOR (15 downto 0);
constant rom : rom_t := (

-- row 0x000
x"0000", x"0000", x"03FC", x"045C", x"0A70", x"0AFC", x"0004", x"0004",
x"0004", x"0004", x"0004", x"0004", x"0104", x"0A74", x"0004", x"0004",

-- row 0x001
x"0004", x"0004", x"0004", x"0004", x"0184", x"0CC4", x"0D44", x"0B44",
x"0B43", x"0C48", x"0337", x"0C44", x"0A1C", x"0AC8", x"008C", x"008C",

-- row 0x002
x"008C", x"008C", x"008C", x"008C", x"008C", x"079C", x"0844", x"08C4",
x"094C", x"03BC", x"0A1C", x"0AC8", x"0088", x"0088", x"0088", x"0088",

-- row 0x003
x"0088", x"0088", x"0088", x"079C", x"0844", x"08C4", x"094C", x"03BC",
x"0A1C", x"0AC8", x"00A0", x"00A0", x"00A0", x"00A0", x"00A0", x"00A0",

-- row 0x004
x"00A0", x"079C", x"0844", x"08C4", x"094C", x"03BC", x"0DC8", x"0A68",
x"0AFC", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0104",

-- row 0x005
x"0A6C", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0184",
x"0B43", x"0B43", x"0337", x"0A08", x"0A8C", x"0788", x"080C", x"08C8",

-- row 0x006
x"0948", x"013C", x"01C0", x"0004", x"0004", x"0004", x"0004", x"0004",
x"0004", x"0984", x"0000", x"0001", x"0A08", x"0A8C", x"0788", x"080C",

-- row 0x007
x"08C8", x"0948", x"013C", x"01C0", x"0005", x"0A08", x"0A8C", x"0788",
x"080C", x"08C8", x"0948", x"013C", x"01C0", x"0004", x"0004", x"0004",

-- row 0x008
x"0004", x"0004", x"0004", x"0484", x"0A08", x"0A8C", x"0788", x"080C",
x"08C8", x"0948", x"013C", x"01C0", x"0004", x"0004", x"0004", x"0004",

-- row 0x009
x"0004", x"0004", x"0504", x"0A24", x"0AA8", x"0005", x"0A08", x"0A8C",
x"0788", x"080C", x"08C8", x"0948", x"013C", x"01C0", x"0004", x"0004",

-- row 0x00A
x"0004", x"0004", x"0004", x"0004", x"0484", x"0A24", x"0AC4", x"0005",
x"0005", x"0005", x"0A08", x"0A8C", x"0788", x"080C", x"08C8", x"0948",

-- row 0x00B
x"013C", x"01C0", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004",
x"0784", x"0844", x"0894", x"0A3C", x"0AC4", x"0004", x"0004", x"0004",

-- row 0x00C
x"0004", x"0004", x"0004", x"0484", x"053C", x"07A8", x"08C8", x"0A3C",
x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0504", x"0A24",

-- row 0x00D
x"0AA8", x"0005", x"0A08", x"0A8C", x"0788", x"080C", x"08C8", x"0948",
x"013C", x"01C0", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004",

-- row 0x00E
x"0484", x"0A24", x"0AC4", x"0004", x"0004", x"0004", x"0004", x"0004",
x"0004", x"0504", x"07A4", x"0844", x"0A3C", x"0004", x"0004", x"0004",

-- row 0x00F
x"0004", x"0004", x"0004", x"0804", x"07A8", x"0898", x"0A3C", x"0AC0",
x"0005", x"0A08", x"0A8C", x"0788", x"080C", x"08C8", x"0948", x"013C",

-- row 0x010
x"01C0", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0784",
x"0894", x"0844", x"0A3C", x"0AC4", x"0005", x"0A08", x"0A8C", x"0788",

-- row 0x011
x"080C", x"08C8", x"0948", x"013C", x"01C0", x"0004", x"0004", x"0004",
x"0004", x"0004", x"0004", x"0484", x"0A08", x"0A8C", x"0788", x"080C",

-- row 0x012
x"08C8", x"0948", x"013C", x"01C0", x"0004", x"0004", x"0004", x"0004",
x"0004", x"0004", x"0504", x"07A4", x"0828", x"0894", x"0A3C", x"0AC0",

-- row 0x013
x"0005", x"0A08", x"0A8C", x"0788", x"080C", x"08C8", x"0948", x"013C",
x"01C0", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0484",

-- row 0x014
x"0A08", x"0A8C", x"0788", x"080C", x"08C8", x"0948", x"013C", x"01C0",
x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0504", x"07A4",

-- row 0x015
x"0828", x"0898", x"0A3C", x"0AC0", x"0005", x"0A08", x"0A8C", x"0788",
x"080C", x"08C8", x"0948", x"013C", x"01C0", x"0004", x"0004", x"0004",

-- row 0x016
x"0004", x"0004", x"0004", x"0884", x"0788", x"080C", x"0D48", x"04BC",
x"0540", x"0D44", x"0005", x"0A08", x"0A8C", x"0788", x"080C", x"08C8",

-- row 0x017
x"0948", x"013C", x"01C0", x"0004", x"0004", x"0004", x"0004", x"0004",
x"0004", x"0484", x"0A08", x"0A8C", x"0788", x"080C", x"08C8", x"0948",

-- row 0x018
x"013C", x"01C0", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004",
x"0504", x"07A4", x"0828", x"08C8", x"0A24", x"0AA8", x"0004", x"0004",

-- row 0x019
x"0004", x"0004", x"0004", x"0004", x"0484", x"0A3C", x"0AC0", x"0004",
x"0004", x"0004", x"0004", x"0004", x"0004", x"0504", x"0A24", x"0AA8",

-- row 0x01A
x"0005", x"0A08", x"0A8C", x"0788", x"080C", x"08C8", x"0948", x"013C",
x"01C0", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0784",

-- row 0x01B
x"0898", x"0844", x"0A3C", x"0AC4", x"0005", x"0004", x"0004", x"0004",
x"0004", x"0004", x"0004", x"0484", x"0009", x"0490", x"0009", x"0790",

-- row 0x01C
x"0844", x"08A4", x"0CA0", x"0948", x"023C", x"05AC", x"0630", x"06B4",
x"0738", x"0CC4", x"000D", x"07A4", x"0890", x"095C", x"023C", x"0630",

-- row 0x01D
x"06B4", x"000D", x"07A4", x"0950", x"04BC", x"05AC", x"0630", x"06B4",
x"000D", x"4047", x"0124", x"01A8", x"000D", x"4046", x"0124", x"01A8",

-- row 0x01E
x"000D", x"404A", x"0124", x"01A8", x"000D", x"07A4", x"0890", x"0958",
x"0630", x"06B4", x"0738", x"000D", x"404E", x"0124", x"01A8", x"000D",

-- row 0x01F
x"404B", x"0124", x"01A8", x"000D", x"404F", x"0124", x"01A8", x"000D",
x"3F03", x"000D", x"4053", x"0124", x"01A8", x"000D", x"4052", x"0124",

-- row 0x020
x"01A8", x"000D", x"000D", x"05C4", x"000D", x"0E44", x"000D", x"0DC4",
x"000D", x"0744", x"000D", x"0790", x"0844", x"08A4", x"0CC8", x"094C",

-- row 0x021
x"05AC", x"0630", x"06B4", x"0CC4", x"000D", x"0794", x"0844", x"08A4",
x"0CC8", x"094C", x"05AC", x"0630", x"06B4", x"0CC4", x"000D", x"0798",

-- row 0x022
x"0844", x"08A4", x"0CC8", x"094C", x"05AC", x"0630", x"06B4", x"0CC4",
x"000D", x"07A4", x"0844", x"08C8", x"0CC8", x"094C", x"04BC", x"0630",

-- row 0x023
x"06B4", x"0CC4", x"000D", x"0794", x"0844", x"08C8", x"0CC8", x"094C",
x"02BC", x"0630", x"06B4", x"0CC4", x"000D", x"0798", x"0844", x"08C8",

-- row 0x024
x"0CC8", x"094C", x"033C", x"0630", x"06B4", x"0CC4", x"000D", x"07A4",
x"0890", x"0964", x"023C", x"0630", x"06B4", x"000D", x"07A4", x"0844",

-- row 0x025
x"08C8", x"0948", x"04BC", x"0630", x"06B4", x"000D", x"0794", x"0844",
x"08C8", x"0948", x"02BC", x"0630", x"06B4", x"000D", x"0798", x"0844",

-- row 0x026
x"08C8", x"0948", x"033C", x"0630", x"06B4", x"000D", x"0124", x"01A8",
x"000D", x"0788", x"080C", x"08C4", x"094C", x"0A1C", x"0AC8", x"00C0",

-- row 0x027
x"00C0", x"00C0", x"00C0", x"00C0", x"00C0", x"00C0", x"079C", x"0844",
x"08C4", x"094C", x"03BC", x"0788", x"080C", x"08C4", x"094C", x"0A1C",

-- row 0x028
x"0AC8", x"00BC", x"00BC", x"00BC", x"00BC", x"00BC", x"00BC", x"00BC",
x"079C", x"0844", x"08C4", x"094C", x"03BC", x"0124", x"01A8", x"000D",

-- row 0x029
x"07A4", x"08C4", x"0948", x"023C", x"0630", x"06B4", x"000D", x"07A4",
x"08C4", x"0948", x"02BC", x"0630", x"06B4", x"000D", x"07A4", x"08C4",

-- row 0x02A
x"0948", x"033C", x"0630", x"06B4", x"000D", x"07A4", x"0954", x"04BC",
x"05AC", x"0630", x"06B4", x"000D", x"000D", x"07A4", x"0890", x"0960",

-- row 0x02B
x"023C", x"0630", x"06B4", x"000D", x"0A1C", x"0AC8", x"079C", x"0844",
x"08C4", x"094C", x"03BC", x"0090", x"0090", x"0090", x"0090", x"0090",

-- row 0x02C
x"0090", x"0090", x"000D", x"0A1C", x"0AC8", x"079C", x"0844", x"08C4",
x"094C", x"03BC", x"00A0", x"00A0", x"00A0", x"00A0", x"00A0", x"00A0",

-- row 0x02D
x"00A0", x"000D", x"079C", x"0844", x"08C8", x"0948", x"03BC", x"0A1C",
x"0AC8", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0784",

-- row 0x02E
x"08C4", x"0948", x"023C", x"0630", x"06B4", x"000D", x"079C", x"0844",
x"08C8", x"0948", x"03BC", x"0A1C", x"0AC8", x"0004", x"0004", x"0004",

-- row 0x02F
x"0004", x"0004", x"0004", x"0404", x"000D", x"07A4", x"0CA0", x"0950",
x"04BC", x"05AC", x"0630", x"06B4", x"0CC4", x"000D", x"07A4", x"0CA0",

-- row 0x030
x"0954", x"04BC", x"05AC", x"0630", x"06B4", x"0CC4", x"000D", x"079C",
x"0844", x"08C8", x"0948", x"03BC", x"0A1C", x"0AC8", x"0004", x"0004",

-- row 0x031
x"0004", x"0004", x"0004", x"0004", x"0404", x"07D8", x"08FC", x"0964",
x"04BC", x"07A0", x"08A4", x"095C", x"043C", x"079C", x"0844", x"08C8",

-- row 0x032
x"0948", x"03BC", x"0A1C", x"0AC8", x"0004", x"0004", x"0004", x"0004",
x"0004", x"0004", x"0104", x"079C", x"0844", x"08C8", x"0948", x"03BC",

-- row 0x033
x"0A1C", x"0AC8", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004",
x"0184", x"000D", x"079C", x"0844", x"08C8", x"0948", x"03BC", x"0A1C",

-- row 0x034
x"0AC8", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0104",
x"079C", x"0844", x"08C8", x"0948", x"03BC", x"0A1C", x"0AC8", x"0004",

-- row 0x035
x"0004", x"0004", x"0004", x"0004", x"0004", x"0184", x"0788", x"080C",
x"08C8", x"0948", x"013C", x"01C0", x"000D", x"0790", x"0844", x"08A4",

-- row 0x036
x"0CA0", x"094C", x"023C", x"05AC", x"0630", x"06B4", x"0738", x"0CC4",
x"000D", x"05C8", x"000D", x"0E48", x"000D", x"0DC8", x"000D", x"0490",

-- row 0x037
x"000D", x"0494", x"000D", x"0498", x"000D", x"0790", x"08C4", x"0948",
x"02BC", x"0630", x"06B4", x"000D", x"0790", x"08C4", x"0948", x"033C",

-- row 0x038
x"0630", x"06B4", x"000D", x"079C", x"08C4", x"0948", x"02BC", x"0630",
x"06B4", x"000D", x"0794", x"08C4", x"0948", x"023C", x"0630", x"06B4",

-- row 0x039
x"000D", x"0394", x"000D", x"0798", x"08C4", x"0948", x"023C", x"0630",
x"06B4", x"000D", x"00A4", x"00A4", x"00A4", x"00A4", x"00A4", x"00A4",

-- row 0x03A
x"00A4", x"0011", x"0224", x"0011", x"0D83", x"36A3", x"37E3", x"0000",
x"0B43", x"0EA3", x"36A3", x"37E3", x"0000", x"0B43", x"12C3", x"36A3",

-- row 0x03B
x"37E3", x"0000", x"0B43", x"1543", x"36A3", x"37E3", x"0000", x"0B43",
x"1A43", x"36A3", x"37E3", x"0000", x"0B43", x"1F23", x"36A3", x"37E3",

-- row 0x03C
x"0000", x"0B43", x"21A3", x"36A3", x"37E3", x"0000", x"0B43", x"2623",
x"36A3", x"37E3", x"0000", x"0B43", x"0D83", x"36A3", x"3963", x"0000",

-- row 0x03D
x"0B43", x"0EA3", x"36A3", x"3963", x"0000", x"0B43", x"12C3", x"36A3",
x"3963", x"0000", x"0B43", x"1543", x"36A3", x"3963", x"0000", x"0B43",

-- row 0x03E
x"1A43", x"36A3", x"3963", x"0000", x"0B43", x"1F23", x"36A3", x"3963",
x"0000", x"0B43", x"21A3", x"36A3", x"3963", x"0000", x"0B43", x"2623",

-- row 0x03F
x"36A3", x"3963", x"0000", x"0B43", x"0EA3", x"36A3", x"3A43", x"7343",
x"0B43", x"12C3", x"36A3", x"3A43", x"7343", x"0B43", x"1503", x"37A3",

-- row 0x040
x"3A43", x"7443", x"0B43", x"1F23", x"36A3", x"3A43", x"7343", x"0B43",
x"21A3", x"36A3", x"3A43", x"7343", x"0B43", x"2AA3", x"0000", x"3B23",

-- row 0x041
x"0000", x"0B43", x"2AA3", x"0000", x"3BA3", x"0000", x"0B43", x"2AA3",
x"0000", x"3C23", x"0000", x"0B43", x"0EA3", x"36A3", x"3CA3", x"0000",

-- row 0x042
x"0B43", x"12C3", x"36A3", x"3CA3", x"0000", x"0B43", x"2AA3", x"0000",
x"3D83", x"0000", x"0B43", x"2AA3", x"0000", x"3E03", x"0000", x"0B43",

-- row 0x043
x"2AA3", x"0000", x"3E83", x"0000", x"0B43", x"1523", x"0000", x"3F03",
x"0000", x"0B43", x"2AA3", x"0000", x"3F43", x"0000", x"0B43", x"2AA3",

-- row 0x044
x"0000", x"3FC3", x"0000", x"0B43", x"1523", x"0000", x"4063", x"0000",
x"0B43", x"1523", x"0000", x"40A3", x"0000", x"0B43", x"1523", x"0000",

-- row 0x045
x"40E3", x"0000", x"0B43", x"1523", x"0000", x"4123", x"0000", x"0B43",
x"0D83", x"36A3", x"4163", x"0000", x"0B43", x"0EA3", x"36A3", x"4163",

-- row 0x046
x"0000", x"0B43", x"12C3", x"36A3", x"4163", x"0000", x"0B43", x"1543",
x"36A3", x"4163", x"0000", x"0B43", x"1A43", x"36A3", x"4163", x"0000",

-- row 0x047
x"0B43", x"1F23", x"36A3", x"4163", x"0000", x"0B43", x"21A3", x"36A3",
x"4163", x"0000", x"0B43", x"2623", x"36A3", x"4163", x"0000", x"0B43",

-- row 0x048
x"0D83", x"36A3", x"42A3", x"0000", x"0B43", x"0EA3", x"36A3", x"42A3",
x"0000", x"0B43", x"12C3", x"36A3", x"42A3", x"0000", x"0B43", x"0D83",

-- row 0x049
x"36A3", x"43E3", x"0000", x"0B43", x"0EA3", x"36A3", x"43E3", x"0000",
x"0B43", x"12C3", x"36A3", x"43E3", x"0000", x"0B43", x"0EA3", x"36A3",

-- row 0x04A
x"4523", x"7343", x"0B43", x"12C3", x"36A3", x"4523", x"7343", x"0B43",
x"1F23", x"36A3", x"4523", x"7343", x"0B43", x"21A3", x"36A3", x"4523",

-- row 0x04B
x"7343", x"0B43", x"1523", x"0000", x"4663", x"0000", x"0B43", x"1523",
x"0000", x"47A3", x"0000", x"0B43", x"0D83", x"36A3", x"48E3", x"0000",

-- row 0x04C
x"0B43", x"0EA3", x"36A3", x"48E3", x"0000", x"0B43", x"12C3", x"36A3",
x"48E3", x"0000", x"0B43", x"1543", x"36A3", x"48E3", x"0000", x"0B43",

-- row 0x04D
x"1A43", x"36A3", x"48E3", x"0000", x"0B43", x"1F23", x"36A3", x"48E3",
x"0000", x"0B43", x"21A3", x"36A3", x"48E3", x"0000", x"0B43", x"2623",

-- row 0x04E
x"36A3", x"48E3", x"0000", x"0B43", x"0EA3", x"36A3", x"49C3", x"7343",
x"0B43", x"12C3", x"36A3", x"49C3", x"7343", x"0B43", x"1F23", x"36A3",

-- row 0x04F
x"49C3", x"7343", x"0B43", x"21A3", x"36A3", x"49C3", x"7343", x"0B43",
x"1523", x"0000", x"4AC3", x"0000", x"0B43", x"1523", x"0000", x"4BC3",

-- row 0x050
x"0000", x"0B43", x"0EA3", x"0000", x"4CC3", x"0000", x"0B43", x"2D63",
x"0000", x"4CC3", x"0000", x"0B43", x"0EA3", x"0000", x"4D23", x"0000",

-- row 0x051
x"0B43", x"0D83", x"36A3", x"5203", x"0000", x"0B43", x"0EA3", x"36A3",
x"5203", x"0000", x"0B43", x"12C3", x"36A3", x"5203", x"0000", x"0B43",

-- row 0x052
x"1543", x"36A3", x"5203", x"0000", x"0B43", x"1A43", x"36A3", x"5203",
x"0000", x"0B43", x"1F23", x"36A3", x"5203", x"0000", x"0B43", x"21A3",

-- row 0x053
x"36A3", x"5203", x"0000", x"0B43", x"2623", x"36A3", x"5203", x"0000",
x"0B43", x"0D83", x"36A3", x"52E3", x"0000", x"0B43", x"0EA3", x"36A3",

-- row 0x054
x"52E3", x"0000", x"0B43", x"12C3", x"36A3", x"52E3", x"0000", x"0B43",
x"2623", x"36A3", x"52E3", x"0000", x"0B43", x"3423", x"36A3", x"52E3",

-- row 0x055
x"0000", x"0B43", x"0D83", x"36A3", x"53C3", x"0000", x"0B43", x"0EA3",
x"36A3", x"53C3", x"0000", x"0B43", x"12C3", x"36A3", x"53C3", x"0000",

-- row 0x056
x"0B43", x"1F23", x"36A3", x"53C3", x"0000", x"0B43", x"21A3", x"36A3",
x"53C3", x"0000", x"0B43", x"0EA3", x"36A3", x"54A3", x"7343", x"0B43",

-- row 0x057
x"12C3", x"36A3", x"54A3", x"7343", x"0B43", x"1503", x"37A3", x"54A3",
x"7443", x"0B43", x"1F23", x"36A3", x"54A3", x"7343", x"0B43", x"21A3",

-- row 0x058
x"36A3", x"54A3", x"7343", x"0B43", x"1523", x"0000", x"5583", x"0000",
x"0B43", x"0D83", x"36A3", x"55A3", x"0000", x"0B43", x"0EA3", x"36A3",

-- row 0x059
x"55A3", x"0000", x"0B43", x"12C3", x"36A3", x"55A3", x"0000", x"0B43",
x"1543", x"36A3", x"55A3", x"0000", x"0B43", x"1A43", x"36A3", x"55A3",

-- row 0x05A
x"0000", x"0B43", x"1F23", x"36A3", x"55A3", x"0000", x"0B43", x"21A3",
x"36A3", x"55A3", x"0000", x"0B43", x"2623", x"36A3", x"55A3", x"0000",

-- row 0x05B
x"0B43", x"1523", x"0000", x"5683", x"0000", x"0B43", x"1523", x"0000",
x"5863", x"0000", x"0B43", x"1523", x"0000", x"5A43", x"0000", x"0B43",

-- row 0x05C
x"1523", x"0000", x"5CC3", x"0000", x"0B43", x"0EA3", x"36A3", x"5EA3",
x"7343", x"0B43", x"12C3", x"36A3", x"5EA3", x"7343", x"0B43", x"1503",

-- row 0x05D
x"37A3", x"5EA3", x"7443", x"0B43", x"1F23", x"36A3", x"5EA3", x"7343",
x"0B43", x"21A3", x"36A3", x"5EA3", x"7343", x"0B43", x"0EA3", x"36A3",

-- row 0x05E
x"5FC3", x"7343", x"0B43", x"12C3", x"36A3", x"5FC3", x"7343", x"0B43",
x"1503", x"37A3", x"5FC3", x"7443", x"0B43", x"1F23", x"36A3", x"5FC3",

-- row 0x05F
x"7343", x"0B43", x"21A3", x"36A3", x"5FC3", x"7343", x"0B43", x"1523",
x"0000", x"60E3", x"0000", x"0B43", x"1523", x"0000", x"6743", x"0000",

-- row 0x060
x"0B43", x"0D83", x"36A3", x"6BA3", x"0000", x"0B43", x"0EA3", x"36A3",
x"6BA3", x"0000", x"0B43", x"12C3", x"36A3", x"6BA3", x"0000", x"0B43",

-- row 0x061
x"1543", x"36A3", x"6BA3", x"0000", x"0B43", x"1A43", x"36A3", x"6BA3",
x"0000", x"0B43", x"1F23", x"36A3", x"6BA3", x"0000", x"0B43", x"21A3",

-- row 0x062
x"36A3", x"6BA3", x"0000", x"0B43", x"2623", x"36A3", x"6BA3", x"0000",
x"0B43", x"1523", x"0000", x"6D23", x"0000", x"0B43", x"1523", x"0000",

-- row 0x063
x"6D63", x"0000", x"0B43", x"1523", x"0000", x"6DA3", x"0000", x"0B43",
x"0EA3", x"0000", x"6DE3", x"7343", x"0B43", x"12C3", x"0000", x"6DE3",

-- row 0x064
x"7343", x"0B43", x"1543", x"0000", x"6DE3", x"7343", x"0B43", x"1A43",
x"0000", x"6DE3", x"7343", x"0B43", x"1F23", x"0000", x"6DE3", x"7343",

-- row 0x065
x"0B43", x"21A3", x"0000", x"6DE3", x"7343", x"0B43", x"2623", x"0000",
x"6DE3", x"7343", x"0B43", x"0EA3", x"0000", x"6E23", x"7343", x"0B43",

-- row 0x066
x"12C3", x"0000", x"6E23", x"7343", x"0B43", x"3423", x"0000", x"6E23",
x"7343", x"0B43", x"0EA3", x"0000", x"6E63", x"7343", x"0B43", x"12C3",

-- row 0x067
x"0000", x"6E63", x"7343", x"0B43", x"1F23", x"0000", x"6E63", x"7343",
x"0B43", x"1523", x"0000", x"6EA3", x"0000", x"0B43", x"1523", x"0000",

-- row 0x068
x"6F83", x"0000", x"0B43", x"1523", x"0000", x"7063", x"0000", x"0B43",
x"1523", x"0000", x"7143", x"0000", x"0B43", x"1523", x"0000", x"7223",

-- row 0x069
x"0000", x"0B43", x"1523", x"0000", x"7263", x"0000", x"0B43", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x06A
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x06B
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x06C
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x06D
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x06E
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x06F
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x070
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x071
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x072
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x073
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x074
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x075
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x076
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x077
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x078
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x079
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x07A
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x07B
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x07C
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x07D
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x07E
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",

-- row 0x07F
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000",
x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000"

);

end package;
