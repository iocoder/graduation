library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

package tlc_test_pkg is
    -- internal signals of vga
    signal VGA_FIRST : STD_LOGIC_VECTOR (7 downto 0);
end package;
