library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

package lookup_pkg is

type rom_t is array (0 to 255) of STD_LOGIC_VECTOR (15 downto 0);
constant rom : rom_t := (

-- row 0x000
x"0435", x"0598", x"0000", x"0000", x"0000", x"0593", x"03F9", x"0000",
x"05B6", x"0589", x"03FE", x"0000", x"0000", x"058E", x"03F4", x"0000",

-- row 0x001
x"0430", x"059D", x"0000", x"0000", x"0000", x"05A2", x"0403", x"0000",
x"0444", x"05AC", x"0000", x"0000", x"0000", x"05A7", x"0408", x"0000",

-- row 0x002
x"050C", x"03DB", x"0000", x"0000", x"0421", x"03D6", x"05CA", x"0000",
x"05C0", x"03CC", x"05CF", x"0000", x"041C", x"03D1", x"05C5", x"0000",

-- row 0x003
x"0426", x"03E0", x"0000", x"0000", x"0000", x"03E5", x"05D4", x"0000",
x"0629", x"03EF", x"0000", x"0000", x"0000", x"03EA", x"05D9", x"0000",

-- row 0x004
x"05F7", x"04CB", x"0000", x"0000", x"0000", x"04C6", x"0570", x"0000",
x"05B1", x"04BC", x"0575", x"0000", x"0502", x"04C1", x"056B", x"0000",

-- row 0x005
x"043A", x"04D0", x"0000", x"0000", x"0000", x"04D5", x"057A", x"0000",
x"044E", x"04DF", x"0000", x"0000", x"0000", x"04DA", x"057F", x"0000",

-- row 0x006
x"05FC", x"03B3", x"0000", x"0000", x"0000", x"03AE", x"05E3", x"0000",
x"05BB", x"03A4", x"05E8", x"0000", x"0507", x"03A9", x"05DE", x"0000",

-- row 0x007
x"043F", x"03B8", x"0000", x"0000", x"0000", x"03BD", x"05ED", x"0000",
x"0633", x"03C7", x"0000", x"0000", x"0000", x"03C2", x"05F2", x"0000",

-- row 0x008
x"0000", x"0642", x"0000", x"0000", x"066F", x"063D", x"0660", x"0000",
x"04B7", x"0000", x"0688", x"0000", x"066A", x"0638", x"065B", x"0000",

-- row 0x009
x"040D", x"0647", x"0000", x"0000", x"0674", x"064C", x"0665", x"0000",
x"0692", x"0656", x"068D", x"0000", x"0000", x"0651", x"0000", x"0000",

-- row 0x00A
x"0552", x"0520", x"0539", x"0000", x"055C", x"051B", x"0543", x"0000",
x"067E", x"0511", x"0679", x"0000", x"0557", x"0516", x"053E", x"0000",

-- row 0x00B
x"0412", x"0525", x"0000", x"0000", x"0561", x"052A", x"054D", x"0000",
x"0453", x"0534", x"0683", x"0000", x"0566", x"052F", x"0548", x"0000",

-- row 0x00C
x"048F", x"0467", x"0000", x"0000", x"0499", x"0462", x"04A3", x"0000",
x"04FD", x"0458", x"04B2", x"0000", x"0494", x"045D", x"049E", x"0000",

-- row 0x00D
x"042B", x"046C", x"0000", x"0000", x"0000", x"0471", x"04A8", x"0000",
x"0449", x"047B", x"0000", x"0000", x"0000", x"0476", x"04AD", x"0000",

-- row 0x00E
x"0480", x"0610", x"0000", x"0000", x"048A", x"060B", x"04E9", x"0000",
x"04F8", x"0601", x"0584", x"0000", x"0485", x"0606", x"04E4", x"0000",

-- row 0x00F
x"0417", x"0615", x"0000", x"0000", x"0000", x"061A", x"04EE", x"0000",
x"062E", x"0624", x"0000", x"0000", x"0000", x"061F", x"04F3", x"0000"

);

end package;
